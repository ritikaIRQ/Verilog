//--------------------------------------------------Hexadecimal to binary encoder------------------------------------------------------------------------------------------------------------------------------

module hex_to_bin(input [15:0] hex,
                  output reg [3:0] bin
                  );

                  always@(*) begin
                    case(hex)
                    16'b0000_0000_0000_0001 : bin = 4'h0;
                    16'b0000_0000_0000_0010 : bin = 4'h1;
                    16'b0000_0000_0000_0100 : bin = 4'h2;
                    16'b0000_0000_0000_1000 : bin = 4'h3;
                    16'b0000_0000_0001_0000 : bin = 4'h4;
                    16'b0000_0000_0010_0000 : bin = 4'h5;
                    16'b0000_0000_0100_0000 : bin = 4'h6;
                    16'b0000_0000_1000_0000 : bin = 4'h7;
                    16'b0000_0001_0000_0000 : bin = 4'h8;
                    16'b0000_0010_0000_0000 : bin = 4'h9;
                    16'b0000_0100_0000_0000 : bin = 4'ha;
                    16'b0000_1000_0000_0000 : bin = 4'hb;
                    16'b0001_0000_0000_0000 : bin = 4'hc;
                    16'b0010_0000_0000_0000 : bin = 4'hd;
                    16'b0100_0000_0000_0000 : bin = 4'he;
                    16'b1000_0000_0000_0000 : bin = 4'hf;
                    default : bin = 4'h0;
                    endcase

                  end

endmodule

