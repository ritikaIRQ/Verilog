//------------------------------------------------------Multiplexer [2:1]-------------------------------------------------------------------------------------------

module mux_2to1(input [1:0] in,
                input sel,
                output y
                );

                assign y = (sel) ? in[1] : in[0];

endmodule